

`include "axis_base_seq.sv"
`include "axis_byte_stream.sv"
`include "axis_cont_aligned_stream.sv"
`include "axis_cont_unaligned_stream.sv"
`include "axis_sparse_stream.sv"