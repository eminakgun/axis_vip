
class axi_cont_unaligned_stream #(`DEFAULT_CLS_PARAM_ARGS) extends axis_base_seq#(`DEFAULT_CLS_PARAMS);
  
  `uvm_object_utils(axis_base_seq#(`DEFAULT_CLS_PARAMS))
  `uvm_object_new

endclass