

`include "axi_base_seq.sv"
`include "axi_byte_stream.sv"
`include "axi_cont_aligned_stream.sv"
`include "axi_cont_unaligned_stream.sv"
`include "axi_sparse_stream.sv"